module preprocess(output wire [3:0] AMod, output wire [3:0] BMod, input wire [3:0] A, input wire [3:0] B, input wire [2:0] Op);

  wire add1;
  wire op1_A;
  wire op2_B,
  wire cpl;

endmodule